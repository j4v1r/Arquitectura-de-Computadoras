----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:56:49 09/30/2025 
-- Design Name: 
-- Module Name:    Ruta - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ruta is
    Port ( clk : in  STD_LOGIC;
           clr : in  STD_LOGIC;
			  s : in STD_LOGIC;
           sd : in  STD_LOGIC_VECTOR (1 downto 0);
           sr : in  STD_LOGIC_VECTOR (1 downto 0);
			  se : in STD_LOGIC_VECTOR (1 downto 0);
           D : in  STD_LOGIC_VECTOR (3 downto 0);
           R : in  STD_LOGIC_VECTOR (3 downto 0);
			  debug_d_aux_antes_suma : out std_logic_vector(3 downto 0);
    debug_r_aux_antes_suma : out std_logic_vector(3 downto 0);
    debug_suma_calculada : out std_logic_vector(4 downto 0);
           N : out  STD_LOGIC;
           C : out  STD_LOGIC;
           Z : out  STD_LOGIC;
           suma : out  STD_LOGIC_VECTOR (3 downto 0));
end ruta;

architecture Behavioral of ruta is

component Registro is
    Port ( clk : in  STD_LOGIC;
           clr : in  STD_LOGIC;
           s1s0 : in  STD_LOGIC_VECTOR (1 downto 0);
           I : in  STD_LOGIC_VECTOR (3 downto 0);
           Q : out  STD_LOGIC_VECTOR (3 downto 0));
end component;

signal Z_aux, N_aux, C_aux : STD_LOGIC;
signal mux_aux, mux_aux_e, d_aux,r_aux, e_aux: std_logic_vector(3 downto 0);
signal suma_aux : std_logic_vector(4 downto 0);

begin

    -- Capturar valores antes de la suma
    process(clk)
    begin
        if rising_edge(clk) then
            if s = '1' then  -- Cuando vamos a hacer suma
                debug_d_aux_antes_suma <= d_aux;
                debug_r_aux_antes_suma <= r_aux;
            end if;
        end if;
    end process;
    
    debug_suma_calculada <= suma_aux;
    
    mux_aux <= D when s='0' else suma_aux(3 downto 0);
    
    suma_aux <= ('0' & d_aux) XOR ('0' & r_aux);
	 
	 Z_aux<=not(suma_aux(3) or suma_aux(2) or suma_aux(1) or suma_aux(0));
	 N_aux<=suma_aux(3);
	 C_aux<=suma_aux(4);
	
	 mux_aux_e<= "0000" when s='0' else ('0'&Z_aux & N_aux & C_aux);
	 
fuente: Registro port map(clk=>clk,clr=>clr,s1s0=>sr,I=>R,Q=>r_aux);
destino: Registro port map(clk=>clk,clr=>clr,s1s0=>sd,I=>mux_aux,Q=>d_aux);
estado: Registro port map(clk=>clk,clr=>clr,s1s0=>se,I=>mux_aux_e,Q=>e_aux);

	Z<=e_aux(2);
	N<=e_aux(1);
	C<=e_aux(0);
	suma<=d_aux;

end Behavioral;

